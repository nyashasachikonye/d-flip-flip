LIBRARY altera;
USE altera.maxplus2.ALL;
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY SCHKUZ_NLSANG001_Lab3_D_Flop IS
	PORT (
		D, CLOCK : IN STD_LOGIC;
		Q, NOTQ : OUT STD_LOGIC
	);
END SCHKUZ_NLSANG001_Lab3_D_Flop;

ARCHITECTURE Behavior OF SCHKUZ_NLSANG001_Lab3_D_Flop IS
BEGIN
	PROCESS (CLOCK)
BEGIN
	IF CLOCK'EVENT AND CLOCK = '1' THEN
		Q <= D;
		NOTQ <= NOT D;
	END IF;
END PROCESS;
END Behavior;
